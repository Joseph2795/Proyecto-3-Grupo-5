`timescale  1 ns / 1 ps
module bcd(clk, number, num);
   // I/O Signal Definitions
   input clk;
   input  [7:0] number;
   output reg [7:0] num;
   
   
always @(posedge clk)  begin
case (number)
8'd0: num <= 8'h00; 
8'd1: num <= 8'h01;
8'd2: num <= 8'h02;
8'd3: num <= 8'h03;
8'd4: num <= 8'h04;
8'd5: num <= 8'h05;
8'd6: num <= 8'h06;
8'd7: num <= 8'h07;
8'd8: num <= 8'h08;
8'd9: num <= 8'h09;
8'd10: num <= 8'h10; 
8'd11: num <= 8'h11;
8'd12: num <= 8'h12;
8'd13: num <= 8'h13;
8'd14: num <= 8'h14;
8'd15: num <= 8'h15;
8'd16: num <= 8'h16;
8'd17: num <= 8'h17;
8'd18: num <= 8'h18;
8'd19: num <= 8'h19;
8'd20: num <= 8'h20; 
8'd21: num <= 8'h21;
8'd22: num <= 8'h22;
8'd23: num <= 8'h23;
8'd24: num <= 8'h24;
8'd25: num <= 8'h25;
8'd26: num <= 8'h26;
8'd27: num <= 8'h27;
8'd28: num <= 8'h28;
8'd29: num <= 8'h29;
8'd30: num <= 8'h30; 
8'd31: num <= 8'h31;
8'd32: num <= 8'h32;
8'd33: num <= 8'h33;
8'd34: num <= 8'h34;
8'd35: num <= 8'h35;
8'd36: num <= 8'h36;
8'd37: num <= 8'h37;
8'd38: num <= 8'h38;
8'd39: num <= 8'h39;
8'd40: num <= 8'h40; 
8'd41: num <= 8'h41;
8'd42: num <= 8'h42;
8'd43: num <= 8'h43;
8'd44: num <= 8'h44;
8'd45: num <= 8'h45;
8'd46: num <= 8'h46;
8'd47: num <= 8'h47;
8'd48: num <= 8'h48;
8'd49: num <= 8'h49;
8'd50: num <= 8'h50; 
8'd51: num <= 8'h51;
8'd52: num <= 8'h52;
8'd53: num <= 8'h53;
8'd54: num <= 8'h54;
8'd55: num <= 8'h55;
8'd56: num <= 8'h56;
8'd57: num <= 8'h57;
8'd58: num <= 8'h58;
8'd59: num <= 8'h59;
8'd60: num <= 8'h60; 
8'd61: num <= 8'h61;
8'd62: num <= 8'h62;
8'd63: num <= 8'h63;
8'd64: num <= 8'h64;
8'd65: num <= 8'h65;
8'd66: num <= 8'h66;
8'd67: num <= 8'h67;
8'd68: num <= 8'h68;
8'd69: num <= 8'h69;
8'd70: num <= 8'h70; 
8'd71: num <= 8'h71;
8'd72: num <= 8'h72;
8'd73: num <= 8'h73;
8'd74: num <= 8'h74;
8'd75: num <= 8'h75;
8'd76: num <= 8'h76;
8'd77: num <= 8'h77;
8'd78: num <= 8'h78;
8'd79: num <= 8'h79;
8'd80: num <= 8'h80; 
8'd81: num <= 8'h81;
8'd82: num <= 8'h82;
8'd83: num <= 8'h83;
8'd84: num <= 8'h84;
8'd85: num <= 8'h85;
8'd86: num <= 8'h86;
8'd87: num <= 8'h87;
8'd88: num <= 8'h88;
8'd89: num <= 8'h89;
8'd90: num <= 8'h90; 
8'd91: num <= 8'h91;
8'd92: num <= 8'h92;
8'd93: num <= 8'h93;
8'd94: num <= 8'h94;
8'd95: num <= 8'h95;
8'd96: num <= 8'h96;
8'd97: num <= 8'h97;
8'd98: num <= 8'h98;
8'd99: num <= 8'h99;
endcase
end
endmodule